module a_gt_eq_six (a2, a1, a0, a_gt_eq_six);
