module something
