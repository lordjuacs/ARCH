module demux16_1x8 (D0,s0,s,y0,y1,y2,y3,y4,y5,y6,y7);
	input[15:0]D0;
	reg [2:0]s;
	output [15:0]y0,y1,y2,y3,y4,y5,y6,y7;

demux	

	F
