module mux16_16x1_not(f,h);
	output f;
	input h;
assign f = ~h;
endmodule
