    Mac OS X            	   2   �      �                                      ATTR       �   �   <                  �   <  com.apple.quarantine q/0083;5ee656ba;Safari;AEAF76F8-01FB-448F-80F4-3DC1B9D06487 