module mux16_8x1_not(f,h);
	output f;
	input h;
assign f = ~h;
endmodule
